module protocol

fn send_ping() {
	
}